*** SPICE deck for cell inv{sch} from library bai_2
*** Created on Thu Oct 23, 2025 20:23:55
*** Last revised on Fri Oct 31, 2025 14:46:33
*** Written on Fri Oct 31, 2025 14:47:05 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inv{sch}
Mnmos-4@0 output input gnd gnd NMOS L=0.6U W=0.6U
Mpmos-4@0 vdd input output vdd PMOS L=0.6U W=1.2U
VDCVoltag@3 vdd gnd DC 5V
VDCVoltag@4 input gnd DC 0V

* Spice Code nodes in cell cell 'inv{sch}'
.op
.include "E:\Analog_IC_Design\ThucHanh\K22_TKVMTT\Electric_2025\libs\models\C5_models.txt"
.END
